class axi_s_wbase_seq extends uvm_sequence #(axi_txn);
  `uvm_object_utils(axi_s_wbase_seq)

  function new(string name = "axi_s_wbase_seq");
    super.new(name);
  endfunction
endclass

